`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07.06.2022 11:04:22
// Design Name: 
// Module Name: Step_input
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Step_input(
    input clk,
    output reg signed [15:0] step_out
    );
    
    /*
    initial begin
        #1;
        step_out = 16'h0000;
    end
    
    initial begin
        #110;
        step_out = 16'hFFEF;
    end
    
    initial begin
        #800;
        step_out = 16'h00FF;
    end
    */
    
    initial begin
        #20;
        step_out = 16'h0080;
        #20;
        step_out = 16'hFF6C;
        #20;
        step_out = 16'h002C;
        #20;
        step_out = 16'h0098;
        #20;
        step_out = 16'h00D9;
        #20;
        step_out = 16'h00BE;
        #20;
        step_out = 16'h004E;
        #20;
        step_out = 16'h018B;
        #20;
        step_out = 16'hFFE7;
        #20;
        step_out = 16'hFFA7;
        #20;
        step_out = 16'h00C5;
        #20;
        step_out = 16'h0038;
        #20;
        step_out = 16'hFF90;
        #20;
        step_out = 16'h0002;
        #20;
        step_out = 16'hFF9E;
        #20;
        step_out = 16'hFFEC;
        #20;
        step_out = 16'h001B;
        #20;
        step_out = 16'h00C5;
        #20;
        step_out = 16'hFFC7;
        #20;
        step_out = 16'h0017;
        #20;
        step_out = 16'h0064;
        #20;
        step_out = 16'hFF44;
        #20;
        step_out = 16'hFF70;
        #20;
        step_out = 16'hFF2A;
        #20;
        step_out = 16'hFFC4;
        #20;
        step_out = 16'hFFE4;
        #20;
        step_out = 16'h004A;
        #20;
        step_out = 16'h0049;
        #20;
        step_out = 16'h00AB;
        #20;
        step_out = 16'h007A;
        #20;
        step_out = 16'hFF2B;
        #20;
        step_out = 16'hFFDC;
        #20;
        step_out = 16'h013C;
        #20;
        step_out = 16'h009F;
        #20;
        step_out = 16'h0099;
        #20;
        step_out = 16'h000F;
        #20;
        step_out = 16'h00DD;
        #20;
        step_out = 16'hFFF6;
        #20;
        step_out = 16'hFFC8;
        #20;
        step_out = 16'hFFCB;
        #20;
        step_out = 16'hFFFA;
        #20;
        step_out = 16'hFF75;
        #20;
        step_out = 16'h009D;
        #20;
        step_out = 16'hFF6C;
        #20;
        step_out = 16'hFEEB;
        #20;
        step_out = 16'hFF1F;
        #20;
        step_out = 16'hFFAB;
        #20;
        step_out = 16'hFF89;
        #20;
        step_out = 16'hFFEE;
        #20;
        step_out = 16'hFF5A;
        #20;
        step_out = 16'hFF8D;
        #20;
        step_out = 16'hFFE1;
        #20;
        step_out = 16'h004A;
        #20;
        step_out = 16'h0021;
        #20;
        step_out = 16'hFFB8;
        #20;
        step_out = 16'h007E;
        #20;
        step_out = 16'hFFEB;
        #20;
        step_out = 16'hFFEC;
        #20;
        step_out = 16'h00CF;
        #20;
        step_out = 16'hFFF2;
        #20;
        step_out = 16'hFF2F;
        #20;
        step_out = 16'hFF9D;
        #20;
        step_out = 16'h0032;
        #20;
        step_out = 16'h001A;
        #20;
        step_out = 16'h0066;
        #20;
        step_out = 16'h00A1;
        #20;
        step_out = 16'h001C;
        #20;
        step_out = 16'h00E5;
        #20;
        step_out = 16'h0016;
        #20;
        step_out = 16'hFFD8;
        #20;
        step_out = 16'h0124;
        #20;
        step_out = 16'h008E;
        #20;
        step_out = 16'h00E2;
        #20;
        step_out = 16'h00BD;
        #20;
        step_out = 16'h007B;
        #20;
        step_out = 16'h0021;
        #20;
        step_out = 16'h009A;
        #20;
        step_out = 16'h00CD;
        #20;
        step_out = 16'h004B;
        #20;
        step_out = 16'h0054;
        #20;
        step_out = 16'h009C;
        #20;
        step_out = 16'h00A0;
        #20;
        step_out = 16'h0030;
        #20;
        step_out = 16'h011E;
        #20;
        step_out = 16'h00A0;
        #20;
        step_out = 16'h0060;
        #20;
        step_out = 16'h0064;
        #20;
        step_out = 16'h0055;
        #20;
        step_out = 16'h002E;
        #20;
        step_out = 16'h0079;
        #20;
        step_out = 16'hFFBF;
        #20;
        step_out = 16'hFFC4;
        #20;
        step_out = 16'hFFEE;
        #20;
        step_out = 16'h0063;
        #20;
        step_out = 16'h004C;
        #20;
        step_out = 16'h00DF;
        #20;
        step_out = 16'h010D;
        #20;
        step_out = 16'h0055;
        #20;
        step_out = 16'hFFB9;
        #20;
        step_out = 16'h0000;
        #20;
        step_out = 16'h0004;
        #20;
        step_out = 16'h0095;
        #20;
        step_out = 16'h0117;
        #20;
        step_out = 16'h00C5;
        #20;
        step_out = 16'h00B3;
        #20;
        step_out = 16'hFF9C;
        #20;
        step_out = 16'hFF5A;
        #20;
        step_out = 16'h008C;
        #20;
        step_out = 16'h00F6;
        #20;
        step_out = 16'hFFB4;
        #20;
        step_out = 16'hFED0;
        #20;
        step_out = 16'hFF8F;
        #20;
        step_out = 16'hFF86;
        #20;
        step_out = 16'hFF39;
        #20;
        step_out = 16'hFFC7;
        #20;
        step_out = 16'h0017;
        #20;
        step_out = 16'hFFBC;
        #20;
        step_out = 16'hFF22;
        #20;
        step_out = 16'hFF8F;
        #20;
        step_out = 16'hFEE2;
        #20;
        step_out = 16'h00D4;
        #20;
        step_out = 16'hFF56;
        #20;
        step_out = 16'h009F;
        #20;
        step_out = 16'hFF87;
        #20;
        step_out = 16'hFFB7;
        #20;
        step_out = 16'hFF82;
        #20;
        step_out = 16'h003D;
        #20;
        step_out = 16'hFF6B;
        #20;
        step_out = 16'hFF73;
        #20;
        step_out = 16'h0008;
        #20;
        step_out = 16'hFFC0;
        #20;
        step_out = 16'h00B7;
        #20;
        step_out = 16'h003F;
        #20;
        step_out = 16'h005C;
        #20;
        step_out = 16'hFF32;
        #20;
        step_out = 16'h0167;
        #20;
        step_out = 16'hFFE2;
        #20;
        step_out = 16'h0074;
        #20;
        step_out = 16'hFFE2;
        #20;
        step_out = 16'h0075;
        #20;
        step_out = 16'hFFB5;
        #20;
        step_out = 16'hFFE1;
        #20;
        step_out = 16'h001C;
        #20;
        step_out = 16'hFF83;
        #20;
        step_out = 16'hFF57;
        #20;
        step_out = 16'h0051;
        #20;
        step_out = 16'h0096;
        #20;
        step_out = 16'hFFBA;
        #20;
        step_out = 16'hFFAB;
        #20;
        step_out = 16'hFFA7;
        #20;
        step_out = 16'hFFC1;
        #20;
        step_out = 16'hFFDB;
        #20;
        step_out = 16'hFF0B;
        #20;
        step_out = 16'hFF64;
        #20;
        step_out = 16'h004F;
        #20;
        step_out = 16'hFFD6;
        #20;
        step_out = 16'hFF4E;
        #20;
        step_out = 16'hFFAB;
        #20;
        step_out = 16'hFFDA;
        #20;
        step_out = 16'h006F;
        #20;
        step_out = 16'h00B9;
        #20;
        step_out = 16'hFF5E;
        #20;
        step_out = 16'hFEEB;
        #20;
        step_out = 16'hFFA8;
        #20;
        step_out = 16'h00A1;
        #20;
        step_out = 16'hFEEA;
        #20;
        step_out = 16'hFF6F;
        #20;
        step_out = 16'h00AC;
        #20;
        step_out = 16'h0049;
        #20;
        step_out = 16'h0005;
        #20;
        step_out = 16'hFFEE;
        #20;
        step_out = 16'h0024;
        #20;
        step_out = 16'h00FE;
        #20;
        step_out = 16'h0016;
        #20;
        step_out = 16'h002F;
        #20;
        step_out = 16'h0055;
        #20;
        step_out = 16'h0133;
        #20;
        step_out = 16'h0014;
        #20;
        step_out = 16'hFF9B;
        #20;
        step_out = 16'h008D;
        #20;
        step_out = 16'hFFD4;
        #20;
        step_out = 16'h0034;
        #20;
        step_out = 16'h001C;
        #20;
        step_out = 16'hFF88;
        #20;
        step_out = 16'h00CC;
        #20;
        step_out = 16'hFFCC;
        #20;
        step_out = 16'h0047;
        #20;
        step_out = 16'hFFFD;
        #20;
        step_out = 16'hFFBC;
        #20;
        step_out = 16'hFFDF;
        #20;
        step_out = 16'h004C;
        #20;
        step_out = 16'h0072;
        #20;
        step_out = 16'hFFA4;
        #20;
        step_out = 16'hFFD8;
        #20;
        step_out = 16'hFFD5;
        #20;
        step_out = 16'h009B;
        #20;
        step_out = 16'h0050;
        #20;
        step_out = 16'h0035;
        #20;
        step_out = 16'h00EA;
        #20;
        step_out = 16'h00C4;
        #20;
        step_out = 16'hFFB4;
        #20;
        step_out = 16'hFF90;
        #20;
        step_out = 16'hFEB4;
        #20;
        step_out = 16'hFF61;
        #20;
        step_out = 16'hFFB5;
        #20;
        step_out = 16'hFFA7;
        #20;
        step_out = 16'h0069;
        #20;
        step_out = 16'hFFA9;
        #20;
        step_out = 16'h0039;
        #20;
        step_out = 16'h0069;
        #20;
        step_out = 16'h0034;
        #20;
        step_out = 16'h0066;
        #20;
        step_out = 16'h011D;
        #20;
        step_out = 16'h0049;
        #20;
        step_out = 16'h00FD;
        #20;
        step_out = 16'h0014;
        #20;
        step_out = 16'hFFC0;
        #20;
        step_out = 16'hFF75;
        #20;
        step_out = 16'hFF00;
        #20;
        step_out = 16'hFFBE;
        #20;
        step_out = 16'h0009;
        #20;
        step_out = 16'hFF9B;
        #20;
        step_out = 16'hFF67;
        #20;
        step_out = 16'h0028;
        #20;
        step_out = 16'h0066;
        #20;
        step_out = 16'hFEC8;
        #20;
        step_out = 16'hFDD2;
        #20;
        step_out = 16'hFF87;
        #20;
        step_out = 16'hFF7B;
        #20;
        step_out = 16'hFF1F;
        #20;
        step_out = 16'h004B;
        #20;
        step_out = 16'h004F;
        #20;
        step_out = 16'hFF74;
        #20;
        step_out = 16'h0051;
        #20;
        step_out = 16'h0065;
        #20;
        step_out = 16'hFFBF;
        #20;
        step_out = 16'hFF5B;
        #20;
        step_out = 16'hFFC3;
        #20;
        step_out = 16'h009A;
        #20;
        step_out = 16'hFFE0;
        #20;
        step_out = 16'hFFC8;
        #20;
        step_out = 16'hFFDA;
        #20;
        step_out = 16'h0069;
        #20;
        step_out = 16'h00B3;
        #20;
        step_out = 16'h0136;
        #20;
        step_out = 16'hFFDC;
        #20;
        step_out = 16'h00DA;
        #20;
        step_out = 16'h0007;
        #20;
        step_out = 16'h003A;
        #20;
        step_out = 16'h0133;
        #20;
        step_out = 16'hFF7B;
        #20;
        step_out = 16'h000D;
        #20;
        step_out = 16'h0074;
        #20;
        step_out = 16'hFF90;
        #20;
        step_out = 16'hFFB9;
        #20;
        step_out = 16'hFF1C;
        #20;
        step_out = 16'h002D;
        #20;
        step_out = 16'hFF52;
        #20;
        step_out = 16'hFED1;
        #20;
        step_out = 16'hFFA0;
        #20;
        step_out = 16'h0045;
        #20;
        step_out = 16'hFF73;
        #20;
        step_out = 16'h0150;
        #20;
        step_out = 16'hFFFE;
        #20;
        step_out = 16'h010B;
        #20;
        step_out = 16'h00B2;
        #20;
        step_out = 16'h010A;
        #20;
        step_out = 16'hFF6F;
        #20;
        step_out = 16'hFF64;
        #20;
        step_out = 16'h00B8;
        #20;
        step_out = 16'hFFBC;
        #20;
        step_out = 16'h00C8;
        #20;
        step_out = 16'h0025;
        #20;
        step_out = 16'hFF68;
        #20;
        step_out = 16'h009A;
        #20;
        step_out = 16'h00DC;
        #20;
        step_out = 16'h0008;
        #20;
        step_out = 16'h012B;
        #20;
        step_out = 16'h00B4;
        #20;
        step_out = 16'hFFD9;
        #20;
        step_out = 16'hFF47;
        #20;
        step_out = 16'hFFF7;
        #20;
        step_out = 16'hFF8C;
        #20;
        step_out = 16'h0163;
        #20;
        step_out = 16'h008C;
        #20;
        step_out = 16'hFF74;
        #20;
        step_out = 16'h0010;
        #20;
        step_out = 16'h01C6;
        #20;
        step_out = 16'h009D;
        #20;
        step_out = 16'h0009;
        #20;
        step_out = 16'hFFF8;
        #20;
        step_out = 16'h0127;
        #20;
        step_out = 16'h00C2;
        #20;
        step_out = 16'h00C8;
        #20;
        step_out = 16'h015D;
        #20;
        step_out = 16'hFFE5;
        #20;
        step_out = 16'h0040;
        #20;
        step_out = 16'h0066;
        #20;
        step_out = 16'h00D0;
        #20;
        step_out = 16'h00C5;
        #20;
        step_out = 16'h0093;
        #20;
        step_out = 16'h009C;
        #20;
        step_out = 16'hFF55;
        #20;
        step_out = 16'hFF29;
        #20;
        step_out = 16'hFE41;
        #20;
        step_out = 16'hFFE7;
        #20;
        step_out = 16'hFF25;
        #20;
        step_out = 16'hFE6D;
        #20;
        step_out = 16'hFFFC;
        #20;
        step_out = 16'h0005;
        #20;
        step_out = 16'h01A0;
        #20;
        step_out = 16'h0118;
        #20;
        step_out = 16'h007C;
        #20;
        step_out = 16'hFFE1;
        #20;
        step_out = 16'hFF65;
        #20;
        step_out = 16'h0043;
        #20;
        step_out = 16'h0047;
        #20;
        step_out = 16'h008E;
        #20;
        step_out = 16'hFF78;
        #20;
        step_out = 16'h007B;
        #20;
        step_out = 16'h00B3;
        #20;
        step_out = 16'h00A2;
        #20;
        step_out = 16'h01B4;
        #20;
        step_out = 16'h0194;
        #20;
        step_out = 16'h00B6;
        #20;
        step_out = 16'h0169;
        #20;
        step_out = 16'h0127;
        #20;
        step_out = 16'h00BB;
        #20;
        step_out = 16'h00AE;
        #20;
        step_out = 16'h0059;
        #20;
        step_out = 16'h0020;
        #20;
        step_out = 16'h0050;
        #20;
        step_out = 16'hFF97;
        #20;
        step_out = 16'hFF4C;
        #20;
        step_out = 16'hFFFF;
        #20;
        step_out = 16'hFF78;
        #20;
        step_out = 16'hFF56;
        #20;
        step_out = 16'h0047;
        #20;
        step_out = 16'hFEF3;
        #20;
        step_out = 16'hFFED;
        #20;
        step_out = 16'hFFD4;
        #20;
        step_out = 16'h00C4;
        #20;
        step_out = 16'h00CD;
        #20;
        step_out = 16'h0195;
        #20;
        step_out = 16'h00D2;
        #20;
        step_out = 16'h011A;
        #20;
        step_out = 16'h0155;
        #20;
        step_out = 16'h00EF;
        #20;
        step_out = 16'h0086;
        #20;
        step_out = 16'h0140;
        #20;
        step_out = 16'h0087;
        #20;
        step_out = 16'h0088;
        #20;
        step_out = 16'h0031;
        #20;
        step_out = 16'h0157;
        #20;
        step_out = 16'h00A6;
        #20;
        step_out = 16'h0091;
        #20;
        step_out = 16'h00B5;
        #20;
        step_out = 16'h0034;
        #20;
        step_out = 16'h00DD;
        #20;
        step_out = 16'h009E;
        #20;
        step_out = 16'hFF34;
        #20;
        step_out = 16'h012B;
        #20;
        step_out = 16'h0141;
        #20;
        step_out = 16'h00B2;
        #20;
        step_out = 16'hFFA5;
        #20;
        step_out = 16'h0049;
        #20;
        step_out = 16'hFFB0;
        #20;
        step_out = 16'h0049;
        #20;
        step_out = 16'hFFD2;
        #20;
        step_out = 16'h0039;
        #20;
        step_out = 16'hFFCE;
        #20;
        step_out = 16'h0054;
        #20;
        step_out = 16'hFFE0;
        #20;
        step_out = 16'hFFA5;
        #20;
        step_out = 16'hFF80;
        #20;
        step_out = 16'hFFC4;
        #20;
        step_out = 16'hFF78;
        #20;
        step_out = 16'h0055;
        #20;
        step_out = 16'h0061;
        #20;
        step_out = 16'h000D;
        #20;
        step_out = 16'h0123;
        #20;
        step_out = 16'h00B9;
        #20;
        step_out = 16'hFFDE;
        #20;
        step_out = 16'hFF5E;
        #20;
        step_out = 16'h00C8;
        #20;
        step_out = 16'h0024;
        #20;
        step_out = 16'hFFD9;
        #20;
        step_out = 16'h0028;
        #20;
        step_out = 16'h008E;
        #20;
        step_out = 16'hFFA9;
        #20;
        step_out = 16'h0026;
        #20;
        step_out = 16'h0051;
        #20;
        step_out = 16'hFEF6;
        #20;
        step_out = 16'hFECA;
        #20;
        step_out = 16'hFF47;
        #20;
        step_out = 16'hFFCA;
        #20;
        step_out = 16'hFF3E;
        #20;
        step_out = 16'h001E;
        #20;
        step_out = 16'h0035;
        #20;
        step_out = 16'hFF7D;
        #20;
        step_out = 16'hFF17;
        #20;
        step_out = 16'h0001;
        #20;
        step_out = 16'hFFE9;
        #20;
        step_out = 16'hFFDD;
        #20;
        step_out = 16'hFE52;
        #20;
        step_out = 16'hFF53;
        #20;
        step_out = 16'hFEF0;
        #20;
        step_out = 16'hFEFE;
        #20;
        step_out = 16'hFFA0;
        #20;
        step_out = 16'h0086;
        #20;
        step_out = 16'hFFD0;
        #20;
        step_out = 16'hFFBE;
        #20;
        step_out = 16'hFFD9;
        #20;
        step_out = 16'h00A2;
        #20;
        step_out = 16'h00D3;
        #20;
        step_out = 16'h0001;
        #20;
        step_out = 16'h012C;
        #20;
        step_out = 16'h0092;
        #20;
        step_out = 16'h00B9;
        #20;
        step_out = 16'h0142;
        #20;
        step_out = 16'hFF19;
        #20;
        step_out = 16'hFF47;
        #20;
        step_out = 16'hFEC7;
        #20;
        step_out = 16'h006E;
        #20;
        step_out = 16'h002D;
        #20;
        step_out = 16'hFFCA;
        #20;
        step_out = 16'h0086;
        #20;
        step_out = 16'hFF70;
        #20;
        step_out = 16'hFEF3;
        #20;
        step_out = 16'hFEFC;
        #20;
        step_out = 16'hFFD1;
        #20;
        step_out = 16'h004F;
        #20;
        step_out = 16'h00EB;
        #20;
        step_out = 16'h007C;
        #20;
        step_out = 16'h0094;
        #20;
        step_out = 16'hFF6A;
        #20;
        step_out = 16'hFE5D;
        #20;
        step_out = 16'hFF9C;
        #20;
        step_out = 16'hFFDF;
        #20;
        step_out = 16'h0044;
        #20;
        step_out = 16'hFF3D;
        #20;
        step_out = 16'h0026;
        #20;
        step_out = 16'h004C;
        #20;
        step_out = 16'h0005;
        #20;
        step_out = 16'h0104;
        #20;
        step_out = 16'h0093;
        #20;
        step_out = 16'h0198;
        #20;
        step_out = 16'h0175;
        #20;
        step_out = 16'hFFC6;
        #20;
        step_out = 16'h00E1;
        #20;
        step_out = 16'h00AA;
        #20;
        step_out = 16'h009F;
        #20;
        step_out = 16'hFF01;
        #20;
        step_out = 16'h001E;
        #20;
        step_out = 16'h0008;
        #20;
        step_out = 16'h0035;
        #20;
        step_out = 16'hFFFF;
        #20;
        step_out = 16'hFFA2;
        #20;
        step_out = 16'h0092;
        #20;
        step_out = 16'hFFD7;
        #20;
        step_out = 16'h009B;
        #20;
        step_out = 16'h002F;
        #20;
        step_out = 16'h0022;
        #20;
        step_out = 16'h0164;
        #20;
        step_out = 16'h00C9;
        #20;
        step_out = 16'h008D;
        #20;
        step_out = 16'h0046;
        #20;
        step_out = 16'h006B;
        #20;
        step_out = 16'hFFDB;
        #20;
        step_out = 16'h0076;
        #20;
        step_out = 16'h004E;
        #20;
        step_out = 16'h013A;
        #20;
        step_out = 16'h0042;
        #20;
        step_out = 16'h0134;
        #20;
        step_out = 16'h003C;
        #20;
        step_out = 16'h00F7;
        #20;
        step_out = 16'hFEE7;
        #20;
        step_out = 16'hFF49;
        #20;
        step_out = 16'hFFBE;
        #20;
        step_out = 16'h0011;
        #20;
        step_out = 16'hFF49;
        #20;
        step_out = 16'h0076;
        #20;
        step_out = 16'h009F;
        #20;
        step_out = 16'hFFEC;
        #20;
        step_out = 16'h005C;
        #20;
        step_out = 16'h00CB;
        #20;
        step_out = 16'h0167;
        #20;
        step_out = 16'h01FA;
        #20;
        step_out = 16'h0119;
        #20;
        step_out = 16'h000F;
        #20;
        step_out = 16'h0060;
        #20;
        step_out = 16'h0047;
        #20;
        step_out = 16'h007C;
        #20;
        step_out = 16'h00A6;
        #20;
        step_out = 16'hFFEC;
        #20;
        step_out = 16'h00BB;
        #20;
        step_out = 16'h0186;
        #20;
        step_out = 16'h00FB;
        #20;
        step_out = 16'h001E;
        #20;
        step_out = 16'h0014;
        #20;
        step_out = 16'hFFB5;
        #20;
        step_out = 16'hFF31;
        #20;
        step_out = 16'hFF23;
        #20;
        step_out = 16'h0059;
        #20;
        step_out = 16'hFFF6;
        #20;
        step_out = 16'h0107;
        #20;
        step_out = 16'hFFD4;
        #20;
        step_out = 16'h0034;
        #20;
        step_out = 16'h004E;
        #20;
        step_out = 16'h020A;
        #20;
        step_out = 16'h015C;
        #20;
        step_out = 16'h00DD;
        #20;
        step_out = 16'h0134;
        #20;
        step_out = 16'h00FD;
        #20;
        step_out = 16'h0138;
        #20;
        step_out = 16'hFFA7;
        #20;
        step_out = 16'hFF9D;
        #20;
        step_out = 16'h009A;
        #20;
        step_out = 16'h00CB;
        #20;
        step_out = 16'h019D;
        #20;
        step_out = 16'hFF8C;
        #20;
        step_out = 16'hFF32;
        #20;
        step_out = 16'hFFD1;
        #20;
        step_out = 16'hFF17;
        #20;
        step_out = 16'h000D;
        #20;
        step_out = 16'h000C;
        #20;
        step_out = 16'hFFFD;
        #20;
        step_out = 16'h006A;
        #20;
        step_out = 16'h004C;
        #20;
        step_out = 16'hFFFC;
        #20;
        step_out = 16'h00FC;
        #20;
        step_out = 16'h007D;
        #20;
        step_out = 16'hFFA5;
        #20;
        step_out = 16'h0015;
        #20;
        step_out = 16'hFFE9;
        #20;
        step_out = 16'h005E;
        #20;
        step_out = 16'hFFC7;
        #20;
        step_out = 16'hFF0C;
        #20;
        step_out = 16'hFF65;
        #20;
        step_out = 16'hFFB8;
        #20;
        step_out = 16'h014D;
        #20;
        step_out = 16'h0022;
        #20;
        step_out = 16'hFFC6;
        #20;
        step_out = 16'hFFED;
        #20;
        step_out = 16'h0040;
        #20;
        step_out = 16'hFFF4;
        #20;
        step_out = 16'h00DE;
        #20;
        step_out = 16'h00AB;
        #20;
        step_out = 16'h01AF;
        #20;
        step_out = 16'h017F;
        #20;
        step_out = 16'h0086;
        #20;
        step_out = 16'h00C8;
        #20;
        step_out = 16'h0062;
        #20;
        step_out = 16'h0015;
        #20;
        step_out = 16'hFFED;
        #20;
        step_out = 16'h018B;
        #20;
        step_out = 16'h006E;
        #20;
        step_out = 16'hFFC9;
        #20;
        step_out = 16'hFFDB;
        #20;
        step_out = 16'h006E;
        #20;
        step_out = 16'h00A1;
        #20;
        step_out = 16'hFFB2;
        #20;
        step_out = 16'hFFEB;
        #20;
        step_out = 16'hFF13;
        #20;
        step_out = 16'h00AB;
        #20;
        step_out = 16'h0005;
        #20;
        step_out = 16'h0025;
        #20;
        step_out = 16'h005E;
        #20;
        step_out = 16'h000F;
        #20;
        step_out = 16'hFF42;
        #20;
        step_out = 16'h001C;
        #20;
        step_out = 16'hFF60;
        #20;
        step_out = 16'h00D1;
        #20;
        step_out = 16'h000F;
        #20;
        step_out = 16'h0142;
        #20;
        step_out = 16'h00F7;
        #20;
        step_out = 16'h0146;
        #20;
        step_out = 16'h0001;
        #20;
        step_out = 16'h0113;
        #20;
        step_out = 16'h0020;
        #20;
        step_out = 16'hFF2A;
        #20;
        step_out = 16'hFFB0;
        #20;
        step_out = 16'h0046;
        #20;
        step_out = 16'hFF58;
        #20;
        step_out = 16'h00CD;
        #20;
        step_out = 16'hFFD0;
        #20;
        step_out = 16'hFFC5;
        #20;
        step_out = 16'hFFDA;
        #20;
        step_out = 16'hFFDF;
        #20;
        step_out = 16'hFF55;
        #20;
        step_out = 16'hFFA5;
        #20;
        step_out = 16'h0062;
        #20;
        step_out = 16'h0012;
        #20;
        step_out = 16'hFFD3;
        #20;
        step_out = 16'h0005;
        #20;
        step_out = 16'h0069;
        #20;
        step_out = 16'h0156;
        #20;
        step_out = 16'h005B;
        #20;
        step_out = 16'h0128;
        #20;
        step_out = 16'h00C5;
        #20;
        step_out = 16'h0013;
        #20;
        step_out = 16'hFFBB;
        #20;
        step_out = 16'h00A2;
        #20;
        step_out = 16'h016F;
        #20;
        step_out = 16'h00CC;
        #20;
        step_out = 16'h009B;
        #20;
        step_out = 16'h00FB;
        #20;
        step_out = 16'h00F6;
        #20;
        step_out = 16'h0069;
        #20;
        step_out = 16'hFF86;
        #20;
        step_out = 16'hFF42;
        #20;
        step_out = 16'h001D;
        #20;
        step_out = 16'hFF8D;
        #20;
        step_out = 16'hFF44;
        #20;
        step_out = 16'hFFB2;
        #20;
        step_out = 16'h000D;
        #20;
        step_out = 16'hFEAF;
        #20;
        step_out = 16'hFF89;
        #20;
        step_out = 16'hFFFA;
        #20;
        step_out = 16'hFF81;
        #20;
        step_out = 16'h00D6;
        #20;
        step_out = 16'h0093;
        #20;
        step_out = 16'h007B;
        #20;
        step_out = 16'h008B;
        #20;
        step_out = 16'hFFFE;
        #20;
        step_out = 16'hFFD8;
        #20;
        step_out = 16'h00FC;
        #20;
        step_out = 16'h0101;
        #20;
        step_out = 16'hFEF0;
        #20;
        step_out = 16'hFF99;
        #20;
        step_out = 16'h001E;
        #20;
        step_out = 16'hFF9E;
        #20;
        step_out = 16'hFFF1;
        #20;
        step_out = 16'h008E;
        #20;
        step_out = 16'h010C;
        #20;
        step_out = 16'h0147;
        #20;
        step_out = 16'h001A;
        #20;
        step_out = 16'h0091;
        #20;
        step_out = 16'h009B;
        #20;
        step_out = 16'h0063;
        #20;
        step_out = 16'h00C3;
        #20;
        step_out = 16'hFFFC;
        #20;
        step_out = 16'h001A;
        #20;
        step_out = 16'hFF74;
        #20;
        step_out = 16'hFFA5;
        #20;
        step_out = 16'h016F;
        #20;
        step_out = 16'h0015;
        #20;
        step_out = 16'h0002;
        #20;
        step_out = 16'hFF81;
        #20;
        step_out = 16'hFF6C;
        #20;
        step_out = 16'hFFEB;
        #20;
        step_out = 16'hFFF6;
        #20;
        step_out = 16'hFFB9;
        #20;
        step_out = 16'hFFC4;
        #20;
        step_out = 16'hFEE7;
        #20;
        step_out = 16'hFF81;
        #20;
        step_out = 16'hFF21;
        #20;
        step_out = 16'hFF13;
        #20;
        step_out = 16'hFFA4;
        #20;
        step_out = 16'hFF24;
        #20;
        step_out = 16'hFF0B;
        #20;
        step_out = 16'h0030;
        #20;
        step_out = 16'hFF8D;
        #20;
        step_out = 16'h00AB;
        #20;
        step_out = 16'hFFB5;
        #20;
        step_out = 16'hFFB9;
        #20;
        step_out = 16'hFE95;
        #20;
        step_out = 16'hFF48;
        #20;
        step_out = 16'hFEF8;
        #20;
        step_out = 16'hFFBB;
        #20;
        step_out = 16'h003E;
        #20;
        step_out = 16'hFFE9;
        #20;
        step_out = 16'hFED5;
        #20;
        step_out = 16'hFF19;
        #20;
        step_out = 16'hFFCD;
        #20;
        step_out = 16'hFEE5;
        #20;
        step_out = 16'hFF64;
        #20;
        step_out = 16'hFEB8;
        #20;
        step_out = 16'hFE92;
        #20;
        step_out = 16'hFF00;
        #20;
        step_out = 16'hFF02;
        #20;
        step_out = 16'hFEEB;
        #20;
        step_out = 16'hFF53;
        #20;
        step_out = 16'hFF44;
        #20;
        step_out = 16'hFEC0;
        #20;
        step_out = 16'hFFA9;
        #20;
        step_out = 16'h007F;
        #20;
        step_out = 16'h006C;
        #20;
        step_out = 16'h002C;
        #20;
        step_out = 16'h0093;
        #20;
        step_out = 16'h0026;
        #20;
        step_out = 16'h015F;
        #20;
        step_out = 16'h002E;
        #20;
        step_out = 16'h0039;
        #20;
        step_out = 16'hFFF4;
        #20;
        step_out = 16'hFFCD;
        #20;
        step_out = 16'h00A4;
        #20;
        step_out = 16'hFFEA;
        #20;
        step_out = 16'hFEE0;
        #20;
        step_out = 16'hFFA9;
        #20;
        step_out = 16'hFF58;
        #20;
        step_out = 16'h006F;
        #20;
        step_out = 16'hFF7C;
        #20;
        step_out = 16'h00DA;
        #20;
        step_out = 16'hFF71;
        #20;
        step_out = 16'hFED2;
        #20;
        step_out = 16'hFF81;
        #20;
        step_out = 16'h0060;
        #20;
        step_out = 16'hFFD2;
        #20;
        step_out = 16'h002D;
        #20;
        step_out = 16'h005C;
        #20;
        step_out = 16'h00A3;
        #20;
        step_out = 16'h008C;
        #20;
        step_out = 16'h0012;
        #20;
        step_out = 16'h000A;
        #20;
        step_out = 16'h0001;
        #20;
        step_out = 16'h0006;
        #20;
        step_out = 16'hFF09;
        #20;
        step_out = 16'hFF48;
        #20;
        step_out = 16'hFEEE;
        #20;
        step_out = 16'h0032;
        #20;
        step_out = 16'hFEB1;
        #20;
        step_out = 16'hFEAE;
        #20;
        step_out = 16'hFF73;
        #20;
        step_out = 16'h0010;
        #20;
        step_out = 16'hFFF9;
        #20;
        step_out = 16'hFFE6;
        #20;
        step_out = 16'hFF1B;
        #20;
        step_out = 16'hFFD0;
        #20;
        step_out = 16'h0022;
        #20;
        step_out = 16'h005B;
        #20;
        step_out = 16'h00DB;
        #20;
        step_out = 16'h003D;
        #20;
        step_out = 16'h0066;
        #20;
        step_out = 16'h0022;
        #20;
        step_out = 16'h006B;
        #20;
        step_out = 16'hFEFD;
        #20;
        step_out = 16'hFF3F;
        #20;
        step_out = 16'h0032;
        #20;
        step_out = 16'h00FA;
        #20;
        step_out = 16'h006B;
        #20;
        step_out = 16'h00B3;
        #20;
        step_out = 16'h001C;
        #20;
        step_out = 16'hFF7C;
        #20;
        step_out = 16'h011E;
        #20;
        step_out = 16'hFFDC;
        #20;
        step_out = 16'hFFDA;
        #20;
        step_out = 16'hFFC7;
        #20;
        step_out = 16'hFFCD;
        #20;
        step_out = 16'hFF8D;
        #20;
        step_out = 16'hFFEF;
        #20;
        step_out = 16'hFF31;
        #20;
        step_out = 16'hFF59;
        #20;
        step_out = 16'hFFA2;
        #20;
        step_out = 16'hFF5F;
        #20;
        step_out = 16'hFF14;
        #20;
        step_out = 16'hFFD8;
        #20;
        step_out = 16'hFEBC;
        #20;
        step_out = 16'hFF6B;
        #20;
        step_out = 16'h006F;
        #20;
        step_out = 16'h0146;
        #20;
        step_out = 16'hFF83;
        #20;
        step_out = 16'h0048;
        #20;
        step_out = 16'h00F0;
        #20;
        step_out = 16'h011E;
        #20;
        step_out = 16'h00B3;
        #20;
        step_out = 16'h0047;
        #20;
        step_out = 16'h001A;
        #20;
        step_out = 16'hFFBE;
        #20;
        step_out = 16'hFF7C;
        #20;
        step_out = 16'hFFC7;
        #20;
        step_out = 16'hFF75;
        #20;
        step_out = 16'h0109;
        #20;
        step_out = 16'h0187;
        #20;
        step_out = 16'h018F;
        #20;
        step_out = 16'h0015;
        #20;
        step_out = 16'hFFFE;
        #20;
        step_out = 16'hFF02;
        #20;
        step_out = 16'hFFFE;
        #20;
        step_out = 16'hFF97;
        #20;
        step_out = 16'h006F;
        #20;
        step_out = 16'h0092;
        #20;
        step_out = 16'hFFAD;
        #20;
        step_out = 16'h006D;
        #20;
        step_out = 16'hFFBB;
        #20;
        step_out = 16'h006E;
        #20;
        step_out = 16'h0161;
        #20;
        step_out = 16'hFFA4;
        #20;
        step_out = 16'h008B;
        #20;
        step_out = 16'h008D;
        #20;
        step_out = 16'h0055;
        #20;
        step_out = 16'h00F4;
        #20;
        step_out = 16'h00D2;
        #20;
        step_out = 16'h0067;
        #20;
        step_out = 16'h00BA;
        #20;
        step_out = 16'hFFE0;
        #20;
        step_out = 16'hFF54;
        #20;
        step_out = 16'hFFEE;
        #20;
        step_out = 16'h0018;
        #20;
        step_out = 16'h0059;
        #20;
        step_out = 16'h007B;
        #20;
        step_out = 16'h00AB;
        #20;
        step_out = 16'h0138;
        #20;
        step_out = 16'h0141;
        #20;
        step_out = 16'h00B1;
        #20;
        step_out = 16'h0053;
        #20;
        step_out = 16'h00AA;
        #20;
        step_out = 16'h0113;
        #20;
        step_out = 16'h0051;
        #20;
        step_out = 16'hFFDE;
        #20;
        step_out = 16'h0002;
        #20;
        step_out = 16'h0069;
        #20;
        step_out = 16'h00AC;
        #20;
        step_out = 16'h00A3;
        #20;
        step_out = 16'h0086;
        #20;
        step_out = 16'hFFF4;
        #20;
        step_out = 16'h0036;
        #20;
        step_out = 16'hFF85;
        #20;
        step_out = 16'hFFE8;
        #20;
        step_out = 16'h009B;
        #20;
        step_out = 16'h01B8;
        #20;
        step_out = 16'h00B0;
        #20;
        step_out = 16'h00C6;
        #20;
        step_out = 16'h00F1;
        #20;
        step_out = 16'h0018;
        #20;
        step_out = 16'h0066;
        #20;
        step_out = 16'h003E;
        #20;
        step_out = 16'h00C9;
        #20;
        step_out = 16'hFF61;
        #20;
        step_out = 16'h00B7;
        #20;
        step_out = 16'h001E;
        #20;
        step_out = 16'hFFCF;
        #20;
        step_out = 16'h00F4;
        #20;
        step_out = 16'h0107;
        #20;
        step_out = 16'h00D0;
        #20;
        step_out = 16'h0147;
        #20;
        step_out = 16'h003F;
        #20;
        step_out = 16'h00B1;
        #20;
        step_out = 16'h00B0;
        #20;
        step_out = 16'h0296;
        #20;
        step_out = 16'h02AE;
        #20;
        step_out = 16'h0198;
        #20;
        step_out = 16'h0264;
        #20;
        step_out = 16'h01C7;
        #20;
        step_out = 16'h00FF;
        #20;
        step_out = 16'h0109;
        #20;
        step_out = 16'h0122;
        #20;
        step_out = 16'h00F4;
        #20;
        step_out = 16'h00E0;
        #20;
        step_out = 16'h00C0;
        #20;
        step_out = 16'h0058;
        #20;
        step_out = 16'h013A;
        #20;
        step_out = 16'h0016;
        #20;
        step_out = 16'h0022;
        #20;
        step_out = 16'h010F;
        #20;
        step_out = 16'h016A;
        #20;
        step_out = 16'h0125;
        #20;
        step_out = 16'h001B;
        #20;
        step_out = 16'h011B;
        #20;
        step_out = 16'h003F;
        #20;
        step_out = 16'hFFFE;
        #20;
        step_out = 16'hFFF4;
        #20;
        step_out = 16'h0033;
        #20;
        step_out = 16'h00D4;
        #20;
        step_out = 16'h0100;
        #20;
        step_out = 16'h002A;
        #20;
        step_out = 16'h007B;
        #20;
        step_out = 16'h002A;
        #20;
        step_out = 16'h006A;
        #20;
        step_out = 16'h009C;
        #20;
        step_out = 16'h002F;
        #20;
        step_out = 16'h00C0;
        #20;
        step_out = 16'h0218;
        #20;
        step_out = 16'h00EF;
        #20;
        step_out = 16'hFF95;
        #20;
        step_out = 16'hFFDB;
        #20;
        step_out = 16'h0097;
        #20;
        step_out = 16'h0015;
        #20;
        step_out = 16'h0067;
        #20;
        step_out = 16'h008E;
        #20;
        step_out = 16'h00BB;
        #20;
        step_out = 16'h0164;
        #20;
        step_out = 16'h005A;
        #20;
        step_out = 16'h010D;
        #20;
        step_out = 16'h012E;
        #20;
        step_out = 16'h01A8;
        #20;
        step_out = 16'h0100;
        #20;
        step_out = 16'h01C6;
        #20;
        step_out = 16'h0077;
        #20;
        step_out = 16'hFFE9;
        #20;
        step_out = 16'h0178;
        #20;
        step_out = 16'h00B8;
        #20;
        step_out = 16'h0030;
        #20;
        step_out = 16'hFFB7;
        #20;
        step_out = 16'hFF20;
        #20;
        step_out = 16'hFFE9;
        #20;
        step_out = 16'h0077;
        #20;
        step_out = 16'h0075;
        #20;
        step_out = 16'h014D;
        #20;
        step_out = 16'h00E5;
        #20;
        step_out = 16'h00FD;
        #20;
        step_out = 16'h014B;
        #20;
        step_out = 16'h0223;
        #20;
        step_out = 16'h012C;
        #20;
        step_out = 16'h0196;
        #20;
        step_out = 16'h016D;
        #20;
        step_out = 16'h0189;
        #20;
        step_out = 16'h023A;
        #20;
        step_out = 16'h00F7;
        #20;
        step_out = 16'h0131;
        #20;
        step_out = 16'h00A8;
        #20;
        step_out = 16'h0001;
        #20;
        step_out = 16'h0033;
        #20;
        step_out = 16'hFF24;
        #20;
        step_out = 16'hFFAE;
        #20;
        step_out = 16'h00D2;
        #20;
        step_out = 16'h003A;
        #20;
        step_out = 16'h0093;
        #20;
        step_out = 16'h0166;
        #20;
        step_out = 16'h01D5;
        #20;
        step_out = 16'h021B;
        #20;
        step_out = 16'h01A7;
        #20;
        step_out = 16'h0185;
        #20;
        step_out = 16'h00ED;
        #20;
        step_out = 16'h0052;
        #20;
        step_out = 16'h0188;
        #20;
        step_out = 16'h0091;
        #20;
        step_out = 16'h015B;
        #20;
        step_out = 16'h01BE;
        #20;
        step_out = 16'h00D8;
        #20;
        step_out = 16'h007D;
        #20;
        step_out = 16'h00A7;
        #20;
        step_out = 16'h00E4;
        #20;
        step_out = 16'h0051;
        #20;
        step_out = 16'h010F;
        #20;
        step_out = 16'h00F2;
        #20;
        step_out = 16'h0108;
        #20;
        step_out = 16'h00A1;
        #20;
        step_out = 16'h00C3;
        #20;
        step_out = 16'h010D;
        #20;
        step_out = 16'h005B;
        #20;
        step_out = 16'h0044;
        #20;
        step_out = 16'h00FC;
        #20;
        step_out = 16'h0071;
        #20;
        step_out = 16'h00C4;
        #20;
        step_out = 16'h0165;
        #20;
        step_out = 16'h0095;
        #20;
        step_out = 16'h00F5;
        #20;
        step_out = 16'h008F;
        #20;
        step_out = 16'h0137;
        #20;
        step_out = 16'h0128;
        #20;
        step_out = 16'h0221;
        #20;
        step_out = 16'h019B;
        #20;
        step_out = 16'h0182;
        #20;
        step_out = 16'h016E;
        #20;
        step_out = 16'h00B8;
        #20;
        step_out = 16'h022D;
        #20;
        step_out = 16'h00EB;
        #20;
        step_out = 16'h0176;
        #20;
        step_out = 16'h0099;
        #20;
        step_out = 16'h00BF;
        #20;
        step_out = 16'h0175;
        #20;
        step_out = 16'h01CA;
        #20;
        step_out = 16'h007F;
        #20;
        step_out = 16'h0176;
        #20;
        step_out = 16'h022A;
        #20;
        step_out = 16'h0186;
        #20;
        step_out = 16'h00F4;
        #20;
        step_out = 16'h00A0;
        #20;
        step_out = 16'h0143;
        #20;
        step_out = 16'h01B7;
        #20;
        step_out = 16'h0105;
        #20;
        step_out = 16'h0151;
        #20;
        step_out = 16'h01CA;
        #20;
        step_out = 16'h017E;
        #20;
        step_out = 16'h01C0;
        #20;
        step_out = 16'h01FE;
        #20;
        step_out = 16'h0149;
        #20;
        step_out = 16'h0270;
        #20;
        step_out = 16'h0259;
        #20;
        step_out = 16'h0140;
        #20;
        step_out = 16'h0131;
        #20;
        step_out = 16'h0266;
        #20;
        step_out = 16'h0173;
        #20;
        step_out = 16'h00EB;
        #20;
        step_out = 16'h0165;
        #20;
        step_out = 16'h014D;
        #20;
        step_out = 16'h0004;
        #20;
        step_out = 16'hFFDA;
        #20;
        step_out = 16'h0075;
        #20;
        step_out = 16'h016A;
        #20;
        step_out = 16'h019F;
        #20;
        step_out = 16'h0176;
        #20;
        step_out = 16'h0161;
        #20;
        step_out = 16'h0239;
        #20;
        step_out = 16'h0125;
        #20;
        step_out = 16'h01DA;
        #20;
        step_out = 16'h011C;
        #20;
        step_out = 16'h01E5;
        #20;
        step_out = 16'h0196;
        #20;
        step_out = 16'h01D3;
        #20;
        step_out = 16'h0260;
        #20;
        step_out = 16'h00A9;
        #20;
        step_out = 16'h02BF;
        #20;
        step_out = 16'h0191;
        #20;
        step_out = 16'h020F;
        #20;
        step_out = 16'h027B;
        #20;
        step_out = 16'h0209;
        #20;
        step_out = 16'h0118;
        #20;
        step_out = 16'h0179;
        #20;
        step_out = 16'h0152;
        #20;
        step_out = 16'h01C8;
        #20;
        step_out = 16'h02AA;
        #20;
        step_out = 16'h0321;
        #20;
        step_out = 16'h02D1;
        #20;
        step_out = 16'h03BE;
        #20;
        step_out = 16'h036C;
        #20;
        step_out = 16'h02FA;
        #20;
        step_out = 16'h03B3;
        #20;
        step_out = 16'h0326;
        #20;
        step_out = 16'h02D1;
        #20;
        step_out = 16'h0370;
        #20;
        step_out = 16'h04A1;
        #20;
        step_out = 16'h0357;
        #20;
        step_out = 16'h03ED;
        #20;
        step_out = 16'h05CF;
        #20;
        step_out = 16'h0548;
        #20;
        step_out = 16'h05AA;
        #20;
        step_out = 16'h074F;
        #20;
        step_out = 16'h0682;
        #20;
        step_out = 16'h078E;
        #20;
        step_out = 16'h07C8;
        #20;
        step_out = 16'h08A8;
        #20;
        step_out = 16'h08D0;
        #20;
        step_out = 16'h096E;
        #20;
        step_out = 16'h08BF;
        #20;
        step_out = 16'h09D2;
        #20;
        step_out = 16'h0BB8;
        #20;
        step_out = 16'h0C28;
        #20;
        step_out = 16'h0BF3;
        #20;
        step_out = 16'h0E33;
        #20;
        step_out = 16'h0D36;
        #20;
        step_out = 16'h0EE6;
        #20;
        step_out = 16'h0EA5;
        #20;
        step_out = 16'h109C;
        #20;
        step_out = 16'h117B;
        #20;
        step_out = 16'h1168;
        #20;
        step_out = 16'h11B1;
        #20;
        step_out = 16'h1163;
        #20;
        step_out = 16'h1217;
        #20;
        step_out = 16'h1299;
        #20;
        step_out = 16'h13D7;
        #20;
        step_out = 16'h12E6;
        #20;
        step_out = 16'h134A;
        #20;
        step_out = 16'h13BF;
        #20;
        step_out = 16'h13F5;
        #20;
        step_out = 16'h13C1;
        #20;
        step_out = 16'h13D7;
        #20;
        step_out = 16'h132E;
        #20;
        step_out = 16'h127D;
        #20;
        step_out = 16'h12F9;
        #20;
        step_out = 16'h12A8;
        #20;
        step_out = 16'h134F;
        #20;
        step_out = 16'h1286;
        #20;
        step_out = 16'h12AD;
        #20;
        step_out = 16'h11DF;
        #20;
        step_out = 16'h124C;
        #20;
        step_out = 16'h1182;
        #20;
        step_out = 16'h1146;
        #20;
        step_out = 16'h103D;
        #20;
        step_out = 16'h0EBA;
        #20;
        step_out = 16'h1003;
        #20;
        step_out = 16'h0EB6;
        #20;
        step_out = 16'h0DB3;
        #20;
        step_out = 16'h0D82;
        #20;
        step_out = 16'h0D3E;
        #20;
        step_out = 16'h0D8B;
        #20;
        step_out = 16'h0DCB;
        #20;
        step_out = 16'h0EF9;
        #20;
        step_out = 16'h0EF5;
        #20;
        step_out = 16'h0E16;
        #20;
        step_out = 16'h0D9B;
        #20;
        step_out = 16'h0DD7;
        #20;
        step_out = 16'h0D65;
        #20;
        step_out = 16'h0D2F;
        #20;
        step_out = 16'h0D94;
        #20;
        step_out = 16'h0D2C;
        #20;
        step_out = 16'h0CB0;
        #20;
        step_out = 16'h0CFB;
        #20;
        step_out = 16'h0BB0;
        #20;
        step_out = 16'h0C66;
        #20;
        step_out = 16'h0C3B;
        #20;
        step_out = 16'h0C32;
        #20;
        step_out = 16'h0C88;
        #20;
        step_out = 16'h0C42;
        #20;
        step_out = 16'h0B80;
        #20;
        step_out = 16'h0B11;
        #20;
        step_out = 16'h0A50;
        #20;
        step_out = 16'h09CE;
        #20;
        step_out = 16'h082F;
        #20;
        step_out = 16'h08FF;
        #20;
        step_out = 16'h0642;
        #20;
        step_out = 16'h0638;
        #20;
        step_out = 16'h0648;
        #20;
        step_out = 16'h064F;
        #20;
        step_out = 16'h063C;
        #20;
        step_out = 16'h054F;
        #20;
        step_out = 16'h0488;
        #20;
        step_out = 16'h0332;
        #20;
        step_out = 16'h02C9;
        #20;
        step_out = 16'h02EC;
        #20;
        step_out = 16'h02C8;
        #20;
        step_out = 16'h02F0;
        #20;
        step_out = 16'h01ED;
        #20;
        step_out = 16'h01EB;
        #20;
        step_out = 16'h0366;
        #20;
        step_out = 16'h02A4;
        #20;
        step_out = 16'h0168;
        #20;
        step_out = 16'h0188;
        #20;
        step_out = 16'h013E;
        #20;
        step_out = 16'h0003;
        #20;
        step_out = 16'hFFBA;
        #20;
        step_out = 16'hFF81;
        #20;
        step_out = 16'hFF4E;
        #20;
        step_out = 16'hFDCA;
        #20;
        step_out = 16'hFD4E;
        #20;
        step_out = 16'hFDEC;
        #20;
        step_out = 16'hFCE4;
        #20;
        step_out = 16'hFD2C;
        #20;
        step_out = 16'hFCA7;
        #20;
        step_out = 16'hFBE1;
        #20;
        step_out = 16'hFB24;
        #20;
        step_out = 16'hFBFB;
        #20;
        step_out = 16'hFA74;
        #20;
        step_out = 16'hFA2B;
        #20;
        step_out = 16'hFB55;
        #20;
        step_out = 16'hFA09;
        #20;
        step_out = 16'hF915;
        #20;
        step_out = 16'hF9D0;
        #20;
        step_out = 16'hFAC4;
        #20;
        step_out = 16'hFA26;
        #20;
        step_out = 16'hF9FB;
        #20;
        step_out = 16'hF9E5;
        #20;
        step_out = 16'hFA09;
        #20;
        step_out = 16'hF98B;
        #20;
        step_out = 16'hF8FF;
        #20;
        step_out = 16'hF9E3;
        #20;
        step_out = 16'hF8E5;
        #20;
        step_out = 16'hF9E3;
        #20;
        step_out = 16'hFA0D;
        #20;
        step_out = 16'hFA07;
        #20;
        step_out = 16'hFA85;
        #20;
        step_out = 16'hF8F5;
        #20;
        step_out = 16'hF998;
        #20;
        step_out = 16'hF9CD;
        #20;
        step_out = 16'hF9B7;
        #20;
        step_out = 16'hFA71;
        #20;
        step_out = 16'hFA6E;
        #20;
        step_out = 16'hFA50;
        #20;
        step_out = 16'hFB6D;
        #20;
        step_out = 16'hFA82;
        #20;
        step_out = 16'hFA0B;
        #20;
        step_out = 16'hFA6D;
        #20;
        step_out = 16'hFB8B;
        #20;
        step_out = 16'hFB70;
        #20;
        step_out = 16'hFAF3;
        #20;
        step_out = 16'hFC1A;
        #20;
        step_out = 16'hFA9D;
        #20;
        step_out = 16'hFAF6;
        #20;
        step_out = 16'hFBF8;
        #20;
        step_out = 16'hFBE3;
        #20;
        step_out = 16'hFC0B;
        #20;
        step_out = 16'hFBF3;
        #20;
        step_out = 16'hFB73;
        #20;
        step_out = 16'hFB5E;
        #20;
        step_out = 16'hFB15;
        #20;
        step_out = 16'hFA9E;
        #20;
        step_out = 16'hFAC7;
        #20;
        step_out = 16'hFAE5;
        #20;
        step_out = 16'hFB1E;
        #20;
        step_out = 16'hFA4D;
        #20;
        step_out = 16'hFA33;
        #20;
        step_out = 16'hFA0F;
        #20;
        step_out = 16'hF9C0;
        #20;
        step_out = 16'hF9D3;
        #20;
        step_out = 16'hF925;
        #20;
        step_out = 16'hF966;
        #20;
        step_out = 16'hF8FC;
        #20;
        step_out = 16'hF9AA;
        #20;
        step_out = 16'hF972;
        #20;
        step_out = 16'hFA5A;
        #20;
        step_out = 16'hFB2D;
        #20;
        step_out = 16'hFA1B;
        #20;
        step_out = 16'hFAE1;
        #20;
        step_out = 16'hFA45;
        #20;
        step_out = 16'hFB27;
        #20;
        step_out = 16'hFAAB;
        #20;
        step_out = 16'hFA68;
        #20;
        step_out = 16'hFA66;
        #20;
        step_out = 16'hFB45;
        #20;
        step_out = 16'hFADB;
        #20;
        step_out = 16'hFB1E;
        #20;
        step_out = 16'hFA17;
        #20;
        step_out = 16'hFA99;
        #20;
        step_out = 16'hF9D3;
        #20;
        step_out = 16'hFA7C;
        #20;
        step_out = 16'hFA59;
        #20;
        step_out = 16'hFA13;
        #20;
        step_out = 16'hFABC;
        #20;
        step_out = 16'hF9E3;
        #20;
        step_out = 16'hF984;
        #20;
        step_out = 16'hFA4A;
        #20;
        step_out = 16'hFB37;
        #20;
        step_out = 16'hF9AF;
        #20;
        step_out = 16'hF96D;
        #20;
        step_out = 16'hF991;
        #20;
        step_out = 16'hFA20;
        #20;
        step_out = 16'hF9AE;
        #20;
        step_out = 16'hF8E0;
        #20;
        step_out = 16'hF92D;
        #20;
        step_out = 16'hFA3F;
        #20;
        step_out = 16'hF9F7;
        #20;
        step_out = 16'hFA1B;
        #20;
        step_out = 16'hF958;
        #20;
        step_out = 16'hF9E8;
        #20;
        step_out = 16'hFAF3;
        #20;
        step_out = 16'hFAC6;
        #20;
        step_out = 16'hFAE9;
        #20;
        step_out = 16'hF87C;
        #20;
        step_out = 16'hF8C2;
        #20;
        step_out = 16'hF945;
        #20;
        step_out = 16'hFA4E;
        #20;
        step_out = 16'hFA5C;
        #20;
        step_out = 16'hF99D;
        #20;
        step_out = 16'hFA80;
        #20;
        step_out = 16'hFACC;
        #20;
        step_out = 16'hFAFA;
        #20;
        step_out = 16'hFA05;
        #20;
        step_out = 16'hF9A3;
        #20;
        step_out = 16'hF9EE;
        #20;
        step_out = 16'hF967;
        #20;
        step_out = 16'hFA94;
        #20;
        step_out = 16'hF8A1;
        #20;
        step_out = 16'hF8CD;
        #20;
        step_out = 16'hF8DB;
        #20;
        step_out = 16'hFA21;
        #20;
        step_out = 16'hF99B;
        #20;
        step_out = 16'hF9B2;
        #20;
        step_out = 16'hF8FF;
        #20;
        step_out = 16'hF992;
        #20;
        step_out = 16'hF916;
        #20;
        step_out = 16'hF964;
        #20;
        step_out = 16'hF887;
        #20;
        step_out = 16'hF85C;
        #20;
        step_out = 16'hF800;
        #20;
        step_out = 16'hF92D;
        #20;
        step_out = 16'hF8D6;
        #20;
        step_out = 16'hF819;
        #20;
        step_out = 16'hF90D;
        #20;
        step_out = 16'hF8D9;
        #20;
        step_out = 16'hF8B3;
        #20;
        step_out = 16'hF7CA;
        #20;
        step_out = 16'hF7E9;
        #20;
        step_out = 16'hF876;
        #20;
        step_out = 16'hF809;
        #20;
        step_out = 16'hF97A;
        #20;
        step_out = 16'hF886;
        #20;
        step_out = 16'hF838;
        #20;
        step_out = 16'hF831;
        #20;
        step_out = 16'hF7FD;
        #20;
        step_out = 16'hF6A0;
        #20;
        step_out = 16'hF788;
        #20;
        step_out = 16'hF79C;
        #20;
        step_out = 16'hF706;
        #20;
        step_out = 16'hF75E;
        #20;
        step_out = 16'hF787;
        #20;
        step_out = 16'hF80B;
        #20;
        step_out = 16'hF82F;
        #20;
        step_out = 16'hF766;
        #20;
        step_out = 16'hF7A1;
        #20;
        step_out = 16'hF7FD;
        #20;
        step_out = 16'hF6D2;
        #20;
        step_out = 16'hF6B0;
        #20;
        step_out = 16'hF76A;
        #20;
        step_out = 16'hF874;
        #20;
        step_out = 16'hF7FB;
        #20;
        step_out = 16'hF91A;
        #20;
        step_out = 16'hF88F;
        #20;
        step_out = 16'hF97A;
        #20;
        step_out = 16'hF78D;
        #20;
        step_out = 16'hF790;
        #20;
        step_out = 16'hF6D5;
        #20;
        step_out = 16'hF747;
        #20;
        step_out = 16'hF70E;
        #20;
        step_out = 16'hF77A;
        #20;
        step_out = 16'hF674;
        #20;
        step_out = 16'hF6F2;
        #20;
        step_out = 16'hF617;
        #20;
        step_out = 16'hF680;
        #20;
        step_out = 16'hF627;
        #20;
        step_out = 16'hF7B0;
        #20;
        step_out = 16'hF74E;
        #20;
        step_out = 16'hF73C;
        #20;
        step_out = 16'hF6D1;
        #20;
        step_out = 16'hF75E;
        #20;
        step_out = 16'hF724;
        #20;
        step_out = 16'hF71D;
        #20;
        step_out = 16'hF76C;
        #20;
        step_out = 16'hF72B;
        #20;
        step_out = 16'hF698;
        #20;
        step_out = 16'hF6A8;
        #20;
        step_out = 16'hF6BD;
        #20;
        step_out = 16'hF701;
        #20;
        step_out = 16'hF701;
        #20;
        step_out = 16'hF5EB;
        #20;
        step_out = 16'hF6C4;
        #20;
        step_out = 16'hF667;
        #20;
        step_out = 16'hF68C;
        #20;
        step_out = 16'hF5FC;
        #20;
        step_out = 16'hF5FF;
        #20;
        step_out = 16'hF721;
        #20;
        step_out = 16'hF7AB;
        #20;
        step_out = 16'hF88A;
        #20;
        step_out = 16'hF880;
        #20;
        step_out = 16'hF789;
        #20;
        step_out = 16'hF7C6;
        #20;
        step_out = 16'hF713;
        #20;
        step_out = 16'hF76E;
        #20;
        step_out = 16'hF6A0;
        #20;
        step_out = 16'hF6FB;
        #20;
        step_out = 16'hF793;
        #20;
        step_out = 16'hF701;
        #20;
        step_out = 16'hF709;
        #20;
        step_out = 16'hF6B4;
        #20;
        step_out = 16'hF70D;
        #20;
        step_out = 16'hF6D2;
        #20;
        step_out = 16'hF576;
        #20;
        step_out = 16'hF6F5;
        #20;
        step_out = 16'hF67A;
        #20;
        step_out = 16'hF65E;
        #20;
        step_out = 16'hF6D8;
        #20;
        step_out = 16'hF674;
        #20;
        step_out = 16'hF53E;
        #20;
        step_out = 16'hF61C;
        #20;
        step_out = 16'hF5E1;
        #20;
        step_out = 16'hF604;
        #20;
        step_out = 16'hF62C;
        #20;
        step_out = 16'hF721;
        #20;
        step_out = 16'hF6A0;
        #20;
        step_out = 16'hF69A;
        #20;
        step_out = 16'hF6D5;
        #20;
        step_out = 16'hF5C6;
        #20;
        step_out = 16'hF5F3;
        #20;
        step_out = 16'hF65B;
        #20;
        step_out = 16'hF6E0;
        #20;
        step_out = 16'hF537;
        #20;
        step_out = 16'hF670;
        #20;
        step_out = 16'hF74C;
        #20;
        step_out = 16'hF504;
        #20;
        step_out = 16'hF5ED;
        #20;
        step_out = 16'hF63C;
        #20;
        step_out = 16'hF6D5;
        #20;
        step_out = 16'hF72E;
        #20;
        step_out = 16'hF64B;
        #20;
        step_out = 16'hF5E7;
        #20;
        step_out = 16'hF612;
        #20;
        step_out = 16'hF5FB;
        #20;
        step_out = 16'hF607;
        #20;
        step_out = 16'hF5C6;
        #20;
        step_out = 16'hF562;
        #20;
        step_out = 16'hF5BA;
        #20;
        step_out = 16'hF61F;
        #20;
        step_out = 16'hF650;
        #20;
        step_out = 16'hF6EB;
        #20;
        step_out = 16'hF69A;
        #20;
        step_out = 16'hF82B;
        #20;
        step_out = 16'hF7AF;
        #20;
        step_out = 16'hF752;
        #20;
        step_out = 16'hF77B;
        #20;
        step_out = 16'hF757;
        #20;
        step_out = 16'hF648;
        #20;
        step_out = 16'hF705;
        #20;
        step_out = 16'hF63C;
        #20;
        step_out = 16'hF72C;
        #20;
        step_out = 16'hF5E3;
        #20;
        step_out = 16'hF648;
        #20;
        step_out = 16'hF6EE;
        #20;
        step_out = 16'hF654;
        #20;
        step_out = 16'hF4D3;
        #20;
        step_out = 16'hF552;
        #20;
        step_out = 16'hF631;
        #20;
        step_out = 16'hF602;
        #20;
        step_out = 16'hF65E;
        #20;
        step_out = 16'hF708;
        #20;
        step_out = 16'hF6BD;
        #20;
        step_out = 16'hF673;
        #20;
        step_out = 16'hF640;
        #20;
        step_out = 16'hF62D;
        #20;
        step_out = 16'hF659;
        #20;
        step_out = 16'hF55F;
        #20;
        step_out = 16'hF4E5;
        #20;
        step_out = 16'hF609;
        #20;
        step_out = 16'hF5EB;
        #20;
        step_out = 16'hF5DA;
        #20;
        step_out = 16'hF5C8;
        #20;
        step_out = 16'hF3FC;
        #20;
        step_out = 16'hF4AC;
        #20;
        step_out = 16'hF5DB;
        #20;
        step_out = 16'hF5DD;
        #20;
        step_out = 16'hF5D4;
        #20;
        step_out = 16'hF5CE;
        #20;
        step_out = 16'hF561;
        #20;
        step_out = 16'hF5B0;
        #20;
        step_out = 16'hF55F;
        #20;
        step_out = 16'hF5C9;
        #20;
        step_out = 16'hF58C;
        #20;
        step_out = 16'hF5A7;
        #20;
        step_out = 16'hF610;
        #20;
        step_out = 16'hF537;
        #20;
        step_out = 16'hF46F;
        #20;
        step_out = 16'hF504;
        #20;
        step_out = 16'hF529;
        #20;
        step_out = 16'hF418;
        #20;
        step_out = 16'hF515;
        #20;
        step_out = 16'hF503;
        #20;
        step_out = 16'hF5F0;
        #20;
        step_out = 16'hF4BE;
        #20;
        step_out = 16'hF454;
        #20;
        step_out = 16'hF383;
        #20;
        step_out = 16'hF4F9;
        #20;
        step_out = 16'hF519;
        #20;
        step_out = 16'hF4CB;
        #20;
        step_out = 16'hF48B;
        #20;
        step_out = 16'hF3F3;
        #20;
        step_out = 16'hF4D0;
        #20;
        step_out = 16'hF4FB;
        #20;
        step_out = 16'hF558;
        #20;
        step_out = 16'hF557;
        #20;
        step_out = 16'hF491;
        #20;
        step_out = 16'hF53B;
        #20;
        step_out = 16'hF48D;
        #20;
        step_out = 16'hF4E2;
        #20;
        step_out = 16'hF442;
        #20;
        step_out = 16'hF661;
        #20;
        step_out = 16'hF5B3;
        #20;
        step_out = 16'hF51A;
        #20;
        step_out = 16'hF5AC;
        #20;
        step_out = 16'hF612;
        #20;
        step_out = 16'hF5EB;
        #20;
        step_out = 16'hF552;
        #20;
        step_out = 16'hF589;
        #20;
        step_out = 16'hF551;
        #20;
        step_out = 16'hF521;
        #20;
        step_out = 16'hF5D4;
        #20;
        step_out = 16'hF52F;
        #20;
        step_out = 16'hF53E;
        #20;
        step_out = 16'hF474;
        #20;
        step_out = 16'hF445;
        #20;
        step_out = 16'hF553;
        #20;
        step_out = 16'hF540;
        #20;
        step_out = 16'hF56F;
        #20;
        step_out = 16'hF5E3;
        #20;
        step_out = 16'hF5E0;
        #20;
        step_out = 16'hF536;
        #20;
        step_out = 16'hF624;
        #20;
        step_out = 16'hF625;
        #20;
        step_out = 16'hF679;
        #20;
        step_out = 16'hF504;
        #20;
        step_out = 16'hF4EF;
        #20;
        step_out = 16'hF4E0;
        #20;
        step_out = 16'hF5A1;
        #20;
        step_out = 16'hF587;
        #20;
        step_out = 16'hF57A;
        #20;
        step_out = 16'hF535;
        #20;
        step_out = 16'hF499;
        #20;
        step_out = 16'hF53E;
        #20;
        step_out = 16'hF527;
        #20;
        step_out = 16'hF4C2;
        #20;
        step_out = 16'hF52A;
        #20;
        step_out = 16'hF530;
        #20;
        step_out = 16'hF544;
        #20;
        step_out = 16'hF49C;
        #20;
        step_out = 16'hF4F5;
        #20;
        step_out = 16'hF49F;
        #20;
        step_out = 16'hF57D;
        #20;
        step_out = 16'hF5EA;
        #20;
        step_out = 16'hF55E;
        #20;
        step_out = 16'hF65D;
        #20;
        step_out = 16'hF514;
        #20;
        step_out = 16'hF5AC;
        #20;
        step_out = 16'hF51E;
        #20;
        step_out = 16'hF447;
        #20;
        step_out = 16'hF481;
        #20;
        step_out = 16'hF404;
        #20;
        step_out = 16'hF557;
        #20;
        step_out = 16'hF3B3;
        #20;
        step_out = 16'hF44D;
        #20;
        step_out = 16'hF440;
        #20;
        step_out = 16'hF3E3;
        #20;
        step_out = 16'hF3FB;
    end
    
endmodule
